module main
import view

fn main() {
	app:=view.new_ui()
	app.run()
}
